// module sshclient
module main // TODO: temporary ...

const (
	version = '0.1.0'
)

fn main() {
	println('Hello World from version $version')
}
